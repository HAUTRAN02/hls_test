// tb.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module tb (
	);

	wire         clock_reset_inst_clock_clk;                                                              // clock_reset_inst:clock -> [component_dpi_controller_pred_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock, mm_host_dpi_bfm_pred_avs_b_conv1_inst:clock, mm_host_dpi_bfm_pred_avs_b_conv2_inst:clock, mm_host_dpi_bfm_pred_avs_b_fc1_inst:clock, mm_host_dpi_bfm_pred_avs_b_fc2_inst:clock, mm_host_dpi_bfm_pred_avs_b_fc3_inst:clock, mm_host_dpi_bfm_pred_avs_image_inst:clock, mm_host_dpi_bfm_pred_avs_probs_inst:clock, mm_host_dpi_bfm_pred_avs_w_conv1_inst:clock, mm_host_dpi_bfm_pred_avs_w_conv2_inst:clock, mm_host_dpi_bfm_pred_avs_w_fc1_inst:clock, mm_host_dpi_bfm_pred_avs_w_fc2_inst:clock, mm_host_dpi_bfm_pred_avs_w_fc3_inst:clock, mm_interconnect_0:clock_reset_inst_clock_clk, mm_interconnect_10:clock_reset_inst_clock_clk, mm_interconnect_11:clock_reset_inst_clock_clk, mm_interconnect_1:clock_reset_inst_clock_clk, mm_interconnect_2:clock_reset_inst_clock_clk, mm_interconnect_3:clock_reset_inst_clock_clk, mm_interconnect_4:clock_reset_inst_clock_clk, mm_interconnect_5:clock_reset_inst_clock_clk, mm_interconnect_6:clock_reset_inst_clock_clk, mm_interconnect_7:clock_reset_inst_clock_clk, mm_interconnect_8:clock_reset_inst_clock_clk, mm_interconnect_9:clock_reset_inst_clock_clk, pred_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                            // clock_reset_inst:clock2x -> [component_dpi_controller_pred_inst:clock2x, main_dpi_controller_inst:clock2x]
	wire         component_dpi_controller_pred_inst_component_call_valid;                                 // component_dpi_controller_pred_inst:start -> pred_inst:start
	wire         pred_inst_call_stall;                                                                    // pred_inst:busy -> component_dpi_controller_pred_inst:busy
	wire         component_dpi_controller_pred_inst_component_done_conduit;                               // component_dpi_controller_pred_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire   [0:0] main_dpi_controller_inst_component_enabled_conduit;                                      // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_pred_inst_component_wait_for_stream_writes_conduit;             // component_dpi_controller_pred_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         component_dpi_controller_pred_inst_dpi_control_bind_conduit;                             // component_dpi_controller_pred_inst:bind_interfaces -> pred_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         mm_host_dpi_bfm_pred_avs_b_conv1_inst_dpi_control_done_reads_conduit;                    // mm_host_dpi_bfm_pred_avs_b_conv1_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_0
	wire         mm_host_dpi_bfm_pred_avs_b_conv2_inst_dpi_control_done_reads_conduit;                    // mm_host_dpi_bfm_pred_avs_b_conv2_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_1
	wire         mm_host_dpi_bfm_pred_avs_w_fc2_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_w_fc2_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_10
	wire         mm_host_dpi_bfm_pred_avs_w_fc3_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_w_fc3_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_11
	wire         mm_host_dpi_bfm_pred_avs_b_fc1_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_b_fc1_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_2
	wire         mm_host_dpi_bfm_pred_avs_b_fc2_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_b_fc2_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_3
	wire         mm_host_dpi_bfm_pred_avs_b_fc3_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_b_fc3_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_4
	wire         mm_host_dpi_bfm_pred_avs_image_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_image_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_5
	wire         mm_host_dpi_bfm_pred_avs_probs_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_probs_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_6
	wire         mm_host_dpi_bfm_pred_avs_w_conv1_inst_dpi_control_done_reads_conduit;                    // mm_host_dpi_bfm_pred_avs_w_conv1_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_7
	wire         mm_host_dpi_bfm_pred_avs_w_conv2_inst_dpi_control_done_reads_conduit;                    // mm_host_dpi_bfm_pred_avs_w_conv2_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_8
	wire         mm_host_dpi_bfm_pred_avs_w_fc1_inst_dpi_control_done_reads_conduit;                      // mm_host_dpi_bfm_pred_avs_w_fc1_inst:done_reads -> pred_component_dpi_controller_agent_done_concatenate_inst:in_conduit_9
	wire         mm_host_dpi_bfm_pred_avs_b_conv1_inst_dpi_control_done_writes_conduit;                   // mm_host_dpi_bfm_pred_avs_b_conv1_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_0
	wire         mm_host_dpi_bfm_pred_avs_b_conv2_inst_dpi_control_done_writes_conduit;                   // mm_host_dpi_bfm_pred_avs_b_conv2_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_1
	wire         mm_host_dpi_bfm_pred_avs_w_fc2_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_w_fc2_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_10
	wire         mm_host_dpi_bfm_pred_avs_w_fc3_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_w_fc3_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_11
	wire         mm_host_dpi_bfm_pred_avs_b_fc1_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_b_fc1_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_2
	wire         mm_host_dpi_bfm_pred_avs_b_fc2_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_b_fc2_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_3
	wire         mm_host_dpi_bfm_pred_avs_b_fc3_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_b_fc3_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_4
	wire         mm_host_dpi_bfm_pred_avs_image_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_image_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_5
	wire         mm_host_dpi_bfm_pred_avs_probs_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_probs_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_6
	wire         mm_host_dpi_bfm_pred_avs_w_conv1_inst_dpi_control_done_writes_conduit;                   // mm_host_dpi_bfm_pred_avs_w_conv1_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_7
	wire         mm_host_dpi_bfm_pred_avs_w_conv2_inst_dpi_control_done_writes_conduit;                   // mm_host_dpi_bfm_pred_avs_w_conv2_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_8
	wire         mm_host_dpi_bfm_pred_avs_w_fc1_inst_dpi_control_done_writes_conduit;                     // mm_host_dpi_bfm_pred_avs_w_fc1_inst:done_writes -> pred_component_dpi_controller_agent_ready_concatenate_inst:in_conduit_9
	wire         component_dpi_controller_pred_inst_dpi_control_enable_conduit;                           // component_dpi_controller_pred_inst:enable_interfaces -> pred_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         concatenate_component_done_inst_out_conduit_conduit;                                     // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire         concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                   // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire  [11:0] pred_component_dpi_controller_agent_done_concatenate_inst_out_conduit_conduit;           // pred_component_dpi_controller_agent_done_concatenate_inst:out_conduit -> component_dpi_controller_pred_inst:agents_done
	wire  [11:0] pred_component_dpi_controller_agent_ready_concatenate_inst_out_conduit_conduit;          // pred_component_dpi_controller_agent_ready_concatenate_inst:out_conduit -> component_dpi_controller_pred_inst:agents_ready
	wire         split_component_start_inst_out_conduit_0_conduit;                                        // split_component_start_inst:out_conduit_0 -> component_dpi_controller_pred_inst:component_enabled
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_0_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_0 -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_1_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_1 -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_10_conduit;           // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_10 -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_10_conduit;         // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_10 -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_10_conduit; // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_10 -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_10_conduit;         // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_10 -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_11_conduit;           // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_11 -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_11_conduit;         // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_11 -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_11_conduit; // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_11 -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_11_conduit;         // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_11 -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_2_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_2 -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_3_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_3 -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_3 -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_4_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_4 -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_4_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_4 -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_5_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_5 -> mm_host_dpi_bfm_pred_avs_image_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_5_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_5 -> mm_host_dpi_bfm_pred_avs_image_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_5_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_5 -> mm_host_dpi_bfm_pred_avs_image_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_5_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_5 -> mm_host_dpi_bfm_pred_avs_image_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_6_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_6 -> mm_host_dpi_bfm_pred_avs_probs_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_6_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_6 -> mm_host_dpi_bfm_pred_avs_probs_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_6_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_6 -> mm_host_dpi_bfm_pred_avs_probs_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_6_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_6 -> mm_host_dpi_bfm_pred_avs_probs_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_7_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_7 -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_7_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_7 -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_7_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_7 -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_7_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_7 -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_8_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_8 -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_8_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_8 -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_8_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_8 -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_8_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_8 -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:enable
	wire         pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_9_conduit;            // pred_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_9 -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:do_bind
	wire         pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_9_conduit;          // pred_component_dpi_controller_agent_readback_fanout_inst:out_conduit_9 -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:component_done
	wire         pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_9_conduit;  // pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_9 -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:component_started
	wire         pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_9_conduit;          // pred_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_9 -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:enable
	wire         component_dpi_controller_pred_inst_read_implicit_streams_conduit;                        // component_dpi_controller_pred_inst:read_implicit_streams -> pred_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_pred_inst_readback_from_agents_conduit;                         // component_dpi_controller_pred_inst:readback_from_agents -> pred_component_dpi_controller_agent_readback_fanout_inst:in_conduit
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                             // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         pred_inst_return_valid;                                                                  // pred_inst:done -> component_dpi_controller_pred_inst:done
	wire         component_dpi_controller_pred_inst_component_return_stall;                               // component_dpi_controller_pred_inst:stall -> pred_inst:stall
	wire         clock_reset_inst_reset_reset;                                                            // clock_reset_inst:resetn -> [component_dpi_controller_pred_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn, mm_host_dpi_bfm_pred_avs_b_conv1_inst:reset_n, mm_host_dpi_bfm_pred_avs_b_conv2_inst:reset_n, mm_host_dpi_bfm_pred_avs_b_fc1_inst:reset_n, mm_host_dpi_bfm_pred_avs_b_fc2_inst:reset_n, mm_host_dpi_bfm_pred_avs_b_fc3_inst:reset_n, mm_host_dpi_bfm_pred_avs_image_inst:reset_n, mm_host_dpi_bfm_pred_avs_probs_inst:reset_n, mm_host_dpi_bfm_pred_avs_w_conv1_inst:reset_n, mm_host_dpi_bfm_pred_avs_w_conv2_inst:reset_n, mm_host_dpi_bfm_pred_avs_w_fc1_inst:reset_n, mm_host_dpi_bfm_pred_avs_w_fc2_inst:reset_n, mm_host_dpi_bfm_pred_avs_w_fc3_inst:reset_n, mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_reset_reset_bridge_in_reset_reset, pred_inst:resetn]
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdata;                                       // mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_waitrequest;                                    // mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_waitrequest
	wire   [4:0] mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_address;                                        // mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_address -> mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_read;                                           // mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_read -> mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_byteenable;                                     // mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_byteenable -> mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdatavalid;                                  // mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_writedata;                                      // mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_writedata -> mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_write;                                          // mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_write -> mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_burstcount;                                     // mm_host_dpi_bfm_pred_avs_b_conv1_inst:avm_burstcount -> mm_interconnect_0:mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_burstcount
	wire  [31:0] mm_interconnect_0_pred_inst_avs_b_conv1_readdata;                                        // pred_inst:avs_b_conv1_readdata -> mm_interconnect_0:pred_inst_avs_b_conv1_readdata
	wire   [2:0] mm_interconnect_0_pred_inst_avs_b_conv1_address;                                         // mm_interconnect_0:pred_inst_avs_b_conv1_address -> pred_inst:avs_b_conv1_address
	wire         mm_interconnect_0_pred_inst_avs_b_conv1_read;                                            // mm_interconnect_0:pred_inst_avs_b_conv1_read -> pred_inst:avs_b_conv1_read
	wire   [3:0] mm_interconnect_0_pred_inst_avs_b_conv1_byteenable;                                      // mm_interconnect_0:pred_inst_avs_b_conv1_byteenable -> pred_inst:avs_b_conv1_byteenable
	wire         mm_interconnect_0_pred_inst_avs_b_conv1_write;                                           // mm_interconnect_0:pred_inst_avs_b_conv1_write -> pred_inst:avs_b_conv1_write
	wire  [31:0] mm_interconnect_0_pred_inst_avs_b_conv1_writedata;                                       // mm_interconnect_0:pred_inst_avs_b_conv1_writedata -> pred_inst:avs_b_conv1_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdata;                                       // mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_waitrequest;                                    // mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_waitrequest
	wire   [5:0] mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_address;                                        // mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_address -> mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_read;                                           // mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_read -> mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_byteenable;                                     // mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_byteenable -> mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdatavalid;                                  // mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_writedata;                                      // mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_writedata -> mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_write;                                          // mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_write -> mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_burstcount;                                     // mm_host_dpi_bfm_pred_avs_b_conv2_inst:avm_burstcount -> mm_interconnect_1:mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_burstcount
	wire  [31:0] mm_interconnect_1_pred_inst_avs_b_conv2_readdata;                                        // pred_inst:avs_b_conv2_readdata -> mm_interconnect_1:pred_inst_avs_b_conv2_readdata
	wire   [3:0] mm_interconnect_1_pred_inst_avs_b_conv2_address;                                         // mm_interconnect_1:pred_inst_avs_b_conv2_address -> pred_inst:avs_b_conv2_address
	wire         mm_interconnect_1_pred_inst_avs_b_conv2_read;                                            // mm_interconnect_1:pred_inst_avs_b_conv2_read -> pred_inst:avs_b_conv2_read
	wire   [3:0] mm_interconnect_1_pred_inst_avs_b_conv2_byteenable;                                      // mm_interconnect_1:pred_inst_avs_b_conv2_byteenable -> pred_inst:avs_b_conv2_byteenable
	wire         mm_interconnect_1_pred_inst_avs_b_conv2_write;                                           // mm_interconnect_1:pred_inst_avs_b_conv2_write -> pred_inst:avs_b_conv2_write
	wire  [31:0] mm_interconnect_1_pred_inst_avs_b_conv2_writedata;                                       // mm_interconnect_1:pred_inst_avs_b_conv2_writedata -> pred_inst:avs_b_conv2_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdata;                                         // mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_waitrequest;                                      // mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_waitrequest
	wire   [8:0] mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_address -> mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_read -> mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_byteenable -> mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdatavalid;                                    // mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_writedata -> mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_write -> mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_b_fc1_inst:avm_burstcount -> mm_interconnect_2:mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_burstcount
	wire  [31:0] mm_interconnect_2_pred_inst_avs_b_fc1_readdata;                                          // pred_inst:avs_b_fc1_readdata -> mm_interconnect_2:pred_inst_avs_b_fc1_readdata
	wire   [6:0] mm_interconnect_2_pred_inst_avs_b_fc1_address;                                           // mm_interconnect_2:pred_inst_avs_b_fc1_address -> pred_inst:avs_b_fc1_address
	wire         mm_interconnect_2_pred_inst_avs_b_fc1_read;                                              // mm_interconnect_2:pred_inst_avs_b_fc1_read -> pred_inst:avs_b_fc1_read
	wire   [3:0] mm_interconnect_2_pred_inst_avs_b_fc1_byteenable;                                        // mm_interconnect_2:pred_inst_avs_b_fc1_byteenable -> pred_inst:avs_b_fc1_byteenable
	wire         mm_interconnect_2_pred_inst_avs_b_fc1_write;                                             // mm_interconnect_2:pred_inst_avs_b_fc1_write -> pred_inst:avs_b_fc1_write
	wire  [31:0] mm_interconnect_2_pred_inst_avs_b_fc1_writedata;                                         // mm_interconnect_2:pred_inst_avs_b_fc1_writedata -> pred_inst:avs_b_fc1_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdata;                                         // mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_waitrequest;                                      // mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_waitrequest
	wire   [8:0] mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_address -> mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_read -> mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_byteenable -> mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdatavalid;                                    // mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_writedata -> mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_write -> mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_b_fc2_inst:avm_burstcount -> mm_interconnect_3:mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_burstcount
	wire  [31:0] mm_interconnect_3_pred_inst_avs_b_fc2_readdata;                                          // pred_inst:avs_b_fc2_readdata -> mm_interconnect_3:pred_inst_avs_b_fc2_readdata
	wire   [6:0] mm_interconnect_3_pred_inst_avs_b_fc2_address;                                           // mm_interconnect_3:pred_inst_avs_b_fc2_address -> pred_inst:avs_b_fc2_address
	wire         mm_interconnect_3_pred_inst_avs_b_fc2_read;                                              // mm_interconnect_3:pred_inst_avs_b_fc2_read -> pred_inst:avs_b_fc2_read
	wire   [3:0] mm_interconnect_3_pred_inst_avs_b_fc2_byteenable;                                        // mm_interconnect_3:pred_inst_avs_b_fc2_byteenable -> pred_inst:avs_b_fc2_byteenable
	wire         mm_interconnect_3_pred_inst_avs_b_fc2_write;                                             // mm_interconnect_3:pred_inst_avs_b_fc2_write -> pred_inst:avs_b_fc2_write
	wire  [31:0] mm_interconnect_3_pred_inst_avs_b_fc2_writedata;                                         // mm_interconnect_3:pred_inst_avs_b_fc2_writedata -> pred_inst:avs_b_fc2_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdata;                                         // mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_waitrequest;                                      // mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_waitrequest
	wire   [5:0] mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_address -> mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_read -> mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_byteenable -> mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdatavalid;                                    // mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_writedata -> mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_write -> mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_b_fc3_inst:avm_burstcount -> mm_interconnect_4:mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_burstcount
	wire  [31:0] mm_interconnect_4_pred_inst_avs_b_fc3_readdata;                                          // pred_inst:avs_b_fc3_readdata -> mm_interconnect_4:pred_inst_avs_b_fc3_readdata
	wire   [3:0] mm_interconnect_4_pred_inst_avs_b_fc3_address;                                           // mm_interconnect_4:pred_inst_avs_b_fc3_address -> pred_inst:avs_b_fc3_address
	wire         mm_interconnect_4_pred_inst_avs_b_fc3_read;                                              // mm_interconnect_4:pred_inst_avs_b_fc3_read -> pred_inst:avs_b_fc3_read
	wire   [3:0] mm_interconnect_4_pred_inst_avs_b_fc3_byteenable;                                        // mm_interconnect_4:pred_inst_avs_b_fc3_byteenable -> pred_inst:avs_b_fc3_byteenable
	wire         mm_interconnect_4_pred_inst_avs_b_fc3_write;                                             // mm_interconnect_4:pred_inst_avs_b_fc3_write -> pred_inst:avs_b_fc3_write
	wire  [31:0] mm_interconnect_4_pred_inst_avs_b_fc3_writedata;                                         // mm_interconnect_4:pred_inst_avs_b_fc3_writedata -> pred_inst:avs_b_fc3_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_image_inst_m0_readdata;                                         // mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_image_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_image_inst_m0_waitrequest;                                      // mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_image_inst:avm_waitrequest
	wire  [11:0] mm_host_dpi_bfm_pred_avs_image_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_image_inst:avm_address -> mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_image_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_image_inst:avm_read -> mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_image_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_image_inst:avm_byteenable -> mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_image_inst_m0_readdatavalid;                                    // mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_image_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_image_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_image_inst:avm_writedata -> mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_image_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_image_inst:avm_write -> mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_image_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_image_inst:avm_burstcount -> mm_interconnect_5:mm_host_dpi_bfm_pred_avs_image_inst_m0_burstcount
	wire  [31:0] mm_interconnect_5_pred_inst_avs_image_readdata;                                          // pred_inst:avs_image_readdata -> mm_interconnect_5:pred_inst_avs_image_readdata
	wire   [9:0] mm_interconnect_5_pred_inst_avs_image_address;                                           // mm_interconnect_5:pred_inst_avs_image_address -> pred_inst:avs_image_address
	wire         mm_interconnect_5_pred_inst_avs_image_read;                                              // mm_interconnect_5:pred_inst_avs_image_read -> pred_inst:avs_image_read
	wire   [3:0] mm_interconnect_5_pred_inst_avs_image_byteenable;                                        // mm_interconnect_5:pred_inst_avs_image_byteenable -> pred_inst:avs_image_byteenable
	wire         mm_interconnect_5_pred_inst_avs_image_write;                                             // mm_interconnect_5:pred_inst_avs_image_write -> pred_inst:avs_image_write
	wire  [31:0] mm_interconnect_5_pred_inst_avs_image_writedata;                                         // mm_interconnect_5:pred_inst_avs_image_writedata -> pred_inst:avs_image_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdata;                                         // mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_probs_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_probs_inst_m0_waitrequest;                                      // mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_probs_inst:avm_waitrequest
	wire   [5:0] mm_host_dpi_bfm_pred_avs_probs_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_probs_inst:avm_address -> mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_probs_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_probs_inst:avm_read -> mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_probs_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_probs_inst:avm_byteenable -> mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdatavalid;                                    // mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_probs_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_probs_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_probs_inst:avm_writedata -> mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_probs_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_probs_inst:avm_write -> mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_probs_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_probs_inst:avm_burstcount -> mm_interconnect_6:mm_host_dpi_bfm_pred_avs_probs_inst_m0_burstcount
	wire  [31:0] mm_interconnect_6_pred_inst_avs_probs_readdata;                                          // pred_inst:avs_probs_readdata -> mm_interconnect_6:pred_inst_avs_probs_readdata
	wire   [3:0] mm_interconnect_6_pred_inst_avs_probs_address;                                           // mm_interconnect_6:pred_inst_avs_probs_address -> pred_inst:avs_probs_address
	wire         mm_interconnect_6_pred_inst_avs_probs_read;                                              // mm_interconnect_6:pred_inst_avs_probs_read -> pred_inst:avs_probs_read
	wire   [3:0] mm_interconnect_6_pred_inst_avs_probs_byteenable;                                        // mm_interconnect_6:pred_inst_avs_probs_byteenable -> pred_inst:avs_probs_byteenable
	wire         mm_interconnect_6_pred_inst_avs_probs_write;                                             // mm_interconnect_6:pred_inst_avs_probs_write -> pred_inst:avs_probs_write
	wire  [31:0] mm_interconnect_6_pred_inst_avs_probs_writedata;                                         // mm_interconnect_6:pred_inst_avs_probs_writedata -> pred_inst:avs_probs_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdata;                                       // mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_waitrequest;                                    // mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_waitrequest
	wire   [4:0] mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_address;                                        // mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_address -> mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_read;                                           // mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_read -> mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_byteenable;                                     // mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_byteenable -> mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdatavalid;                                  // mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_writedata;                                      // mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_writedata -> mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_write;                                          // mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_write -> mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_burstcount;                                     // mm_host_dpi_bfm_pred_avs_w_conv1_inst:avm_burstcount -> mm_interconnect_7:mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_burstcount
	wire  [31:0] mm_interconnect_7_pred_inst_avs_w_conv1_readdata;                                        // pred_inst:avs_w_conv1_readdata -> mm_interconnect_7:pred_inst_avs_w_conv1_readdata
	wire   [2:0] mm_interconnect_7_pred_inst_avs_w_conv1_address;                                         // mm_interconnect_7:pred_inst_avs_w_conv1_address -> pred_inst:avs_w_conv1_address
	wire         mm_interconnect_7_pred_inst_avs_w_conv1_read;                                            // mm_interconnect_7:pred_inst_avs_w_conv1_read -> pred_inst:avs_w_conv1_read
	wire   [3:0] mm_interconnect_7_pred_inst_avs_w_conv1_byteenable;                                      // mm_interconnect_7:pred_inst_avs_w_conv1_byteenable -> pred_inst:avs_w_conv1_byteenable
	wire         mm_interconnect_7_pred_inst_avs_w_conv1_write;                                           // mm_interconnect_7:pred_inst_avs_w_conv1_write -> pred_inst:avs_w_conv1_write
	wire  [31:0] mm_interconnect_7_pred_inst_avs_w_conv1_writedata;                                       // mm_interconnect_7:pred_inst_avs_w_conv1_writedata -> pred_inst:avs_w_conv1_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdata;                                       // mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_waitrequest;                                    // mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_waitrequest
	wire  [13:0] mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_address;                                        // mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_address -> mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_read;                                           // mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_read -> mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_byteenable;                                     // mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_byteenable -> mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdatavalid;                                  // mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_writedata;                                      // mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_writedata -> mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_write;                                          // mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_write -> mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_burstcount;                                     // mm_host_dpi_bfm_pred_avs_w_conv2_inst:avm_burstcount -> mm_interconnect_8:mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_burstcount
	wire  [31:0] mm_interconnect_8_pred_inst_avs_w_conv2_readdata;                                        // pred_inst:avs_w_conv2_readdata -> mm_interconnect_8:pred_inst_avs_w_conv2_readdata
	wire  [11:0] mm_interconnect_8_pred_inst_avs_w_conv2_address;                                         // mm_interconnect_8:pred_inst_avs_w_conv2_address -> pred_inst:avs_w_conv2_address
	wire         mm_interconnect_8_pred_inst_avs_w_conv2_read;                                            // mm_interconnect_8:pred_inst_avs_w_conv2_read -> pred_inst:avs_w_conv2_read
	wire   [3:0] mm_interconnect_8_pred_inst_avs_w_conv2_byteenable;                                      // mm_interconnect_8:pred_inst_avs_w_conv2_byteenable -> pred_inst:avs_w_conv2_byteenable
	wire         mm_interconnect_8_pred_inst_avs_w_conv2_write;                                           // mm_interconnect_8:pred_inst_avs_w_conv2_write -> pred_inst:avs_w_conv2_write
	wire  [31:0] mm_interconnect_8_pred_inst_avs_w_conv2_writedata;                                       // mm_interconnect_8:pred_inst_avs_w_conv2_writedata -> pred_inst:avs_w_conv2_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdata;                                         // mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_waitrequest;                                      // mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_waitrequest
	wire  [17:0] mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_address -> mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_read -> mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_byteenable -> mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdatavalid;                                    // mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_writedata -> mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_write -> mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_w_fc1_inst:avm_burstcount -> mm_interconnect_9:mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_burstcount
	wire  [31:0] mm_interconnect_9_pred_inst_avs_w_fc1_readdata;                                          // pred_inst:avs_w_fc1_readdata -> mm_interconnect_9:pred_inst_avs_w_fc1_readdata
	wire  [15:0] mm_interconnect_9_pred_inst_avs_w_fc1_address;                                           // mm_interconnect_9:pred_inst_avs_w_fc1_address -> pred_inst:avs_w_fc1_address
	wire         mm_interconnect_9_pred_inst_avs_w_fc1_read;                                              // mm_interconnect_9:pred_inst_avs_w_fc1_read -> pred_inst:avs_w_fc1_read
	wire   [3:0] mm_interconnect_9_pred_inst_avs_w_fc1_byteenable;                                        // mm_interconnect_9:pred_inst_avs_w_fc1_byteenable -> pred_inst:avs_w_fc1_byteenable
	wire         mm_interconnect_9_pred_inst_avs_w_fc1_write;                                             // mm_interconnect_9:pred_inst_avs_w_fc1_write -> pred_inst:avs_w_fc1_write
	wire  [31:0] mm_interconnect_9_pred_inst_avs_w_fc1_writedata;                                         // mm_interconnect_9:pred_inst_avs_w_fc1_writedata -> pred_inst:avs_w_fc1_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdata;                                         // mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_waitrequest;                                      // mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_waitrequest
	wire  [15:0] mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_address -> mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_read -> mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_byteenable -> mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdatavalid;                                    // mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_writedata -> mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_write -> mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_w_fc2_inst:avm_burstcount -> mm_interconnect_10:mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_burstcount
	wire  [31:0] mm_interconnect_10_pred_inst_avs_w_fc2_readdata;                                         // pred_inst:avs_w_fc2_readdata -> mm_interconnect_10:pred_inst_avs_w_fc2_readdata
	wire  [13:0] mm_interconnect_10_pred_inst_avs_w_fc2_address;                                          // mm_interconnect_10:pred_inst_avs_w_fc2_address -> pred_inst:avs_w_fc2_address
	wire         mm_interconnect_10_pred_inst_avs_w_fc2_read;                                             // mm_interconnect_10:pred_inst_avs_w_fc2_read -> pred_inst:avs_w_fc2_read
	wire   [3:0] mm_interconnect_10_pred_inst_avs_w_fc2_byteenable;                                       // mm_interconnect_10:pred_inst_avs_w_fc2_byteenable -> pred_inst:avs_w_fc2_byteenable
	wire         mm_interconnect_10_pred_inst_avs_w_fc2_write;                                            // mm_interconnect_10:pred_inst_avs_w_fc2_write -> pred_inst:avs_w_fc2_write
	wire  [31:0] mm_interconnect_10_pred_inst_avs_w_fc2_writedata;                                        // mm_interconnect_10:pred_inst_avs_w_fc2_writedata -> pred_inst:avs_w_fc2_writedata
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdata;                                         // mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdata -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_readdata
	wire         mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_waitrequest;                                      // mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_waitrequest -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_waitrequest
	wire  [11:0] mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_address;                                          // mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_address -> mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_address
	wire         mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_read;                                             // mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_read -> mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_read
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_byteenable;                                       // mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_byteenable -> mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_byteenable
	wire         mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdatavalid;                                    // mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdatavalid -> mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_readdatavalid
	wire   [7:0] mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_writedata;                                        // mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_writedata -> mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_writedata
	wire         mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_write;                                            // mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_write -> mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_write
	wire   [0:0] mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_burstcount;                                       // mm_host_dpi_bfm_pred_avs_w_fc3_inst:avm_burstcount -> mm_interconnect_11:mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_burstcount
	wire  [31:0] mm_interconnect_11_pred_inst_avs_w_fc3_readdata;                                         // pred_inst:avs_w_fc3_readdata -> mm_interconnect_11:pred_inst_avs_w_fc3_readdata
	wire   [9:0] mm_interconnect_11_pred_inst_avs_w_fc3_address;                                          // mm_interconnect_11:pred_inst_avs_w_fc3_address -> pred_inst:avs_w_fc3_address
	wire         mm_interconnect_11_pred_inst_avs_w_fc3_read;                                             // mm_interconnect_11:pred_inst_avs_w_fc3_read -> pred_inst:avs_w_fc3_read
	wire   [3:0] mm_interconnect_11_pred_inst_avs_w_fc3_byteenable;                                       // mm_interconnect_11:pred_inst_avs_w_fc3_byteenable -> pred_inst:avs_w_fc3_byteenable
	wire         mm_interconnect_11_pred_inst_avs_w_fc3_write;                                            // mm_interconnect_11:pred_inst_avs_w_fc3_write -> pred_inst:avs_w_fc3_write
	wire  [31:0] mm_interconnect_11_pred_inst_avs_w_fc3_writedata;                                        // mm_interconnect_11:pred_inst_avs_w_fc3_writedata -> pred_inst:avs_w_fc3_writedata
	wire         component_dpi_controller_pred_inst_component_irq_irq;                                    // irq_mapper:sender_irq -> component_dpi_controller_pred_inst:done_irq

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("pred"),
		.COMPONENT_MANGLED_NAME       ("\\3fpred@@YAXPEAM00000000000@Z"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (12),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_pred_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                     //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                   //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                   //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_pred_inst_dpi_control_bind_conduit),                    //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_pred_inst_dpi_control_enable_conduit),                  //               dpi_control_enable.conduit
		.agents_ready                     (pred_component_dpi_controller_agent_ready_concatenate_inst_out_conduit_conduit), //         dpi_control_agents_ready.conduit
		.agents_done                      (pred_component_dpi_controller_agent_done_concatenate_inst_out_conduit_conduit),  //          dpi_control_agents_done.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                               //                component_enabled.conduit
		.component_done                   (component_dpi_controller_pred_inst_component_done_conduit),                      //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_pred_inst_component_wait_for_stream_writes_conduit),    // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                               //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_pred_inst_read_implicit_streams_conduit),               //            read_implicit_streams.conduit
		.readback_from_agents             (component_dpi_controller_pred_inst_readback_from_agents_conduit),                //             readback_from_agents.conduit
		.start                            (component_dpi_controller_pred_inst_component_call_valid),                        //                   component_call.valid
		.busy                             (pred_inst_call_stall),                                                           //                                 .stall
		.done                             (pred_inst_return_valid),                                                         //                 component_return.valid
		.stall                            (component_dpi_controller_pred_inst_component_return_stall),                      //                                 .stall
		.done_irq                         (component_dpi_controller_pred_inst_component_irq_irq),                           //                    component_irq.irq
		.returndata                       ()                                                                                //                       returndata.data
	);

	tb_concatenate_component_done_inst concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),       //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_pred_inst_component_done_conduit)  // in_conduit_0.conduit
	);

	tb_concatenate_component_done_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),       //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_pred_inst_component_wait_for_stream_writes_conduit)  // in_conduit_0.conduit
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS      (1),
		.COMPONENT_NAMES_STR ("pred")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (5),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("b_conv1"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("b_conv1_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_b_conv1_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_b_conv1_inst_dpi_control_done_writes_conduit),                  //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_b_conv1_inst_dpi_control_done_reads_conduit),                   //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_0_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_writedata),                                     //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_burstcount),                                    //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdata),                                      //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_address),                                       //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_waitrequest),                                   //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_write),                                         //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_read),                                          //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_byteenable),                                    //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdatavalid)                                  //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (6),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("b_conv2"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("b_conv2_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_b_conv2_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_b_conv2_inst_dpi_control_done_writes_conduit),                  //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_b_conv2_inst_dpi_control_done_reads_conduit),                   //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_1_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_writedata),                                     //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_burstcount),                                    //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdata),                                      //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_address),                                       //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_waitrequest),                                   //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_write),                                         //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_read),                                          //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_byteenable),                                    //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdatavalid)                                  //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (9),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("b_fc1"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("b_fc1_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_b_fc1_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_b_fc1_inst_dpi_control_done_writes_conduit),                    //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_b_fc1_inst_dpi_control_done_reads_conduit),                     //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_2_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_writedata),                                       //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_burstcount),                                      //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdata),                                        //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_address),                                         //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_waitrequest),                                     //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_write),                                           //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_read),                                            //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_byteenable),                                      //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdatavalid)                                    //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (9),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("b_fc2"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("b_fc2_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_b_fc2_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_b_fc2_inst_dpi_control_done_writes_conduit),                    //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_b_fc2_inst_dpi_control_done_reads_conduit),                     //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_3_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_writedata),                                       //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_burstcount),                                      //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdata),                                        //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_address),                                         //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_waitrequest),                                     //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_write),                                           //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_read),                                            //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_byteenable),                                      //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdatavalid)                                    //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (6),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("b_fc3"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("b_fc3_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_b_fc3_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_b_fc3_inst_dpi_control_done_writes_conduit),                    //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_b_fc3_inst_dpi_control_done_reads_conduit),                     //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_4_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_4_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_writedata),                                       //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_burstcount),                                      //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdata),                                        //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_address),                                         //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_waitrequest),                                     //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_write),                                           //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_read),                                            //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_byteenable),                                      //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdatavalid)                                    //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (12),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("image"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("image_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_image_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_5_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_5_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_image_inst_dpi_control_done_writes_conduit),                    //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_image_inst_dpi_control_done_reads_conduit),                     //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_5_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_5_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_image_inst_m0_writedata),                                       //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_image_inst_m0_burstcount),                                      //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_image_inst_m0_readdata),                                        //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_image_inst_m0_address),                                         //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_image_inst_m0_waitrequest),                                     //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_image_inst_m0_write),                                           //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_image_inst_m0_read),                                            //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_image_inst_m0_byteenable),                                      //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_image_inst_m0_readdatavalid)                                    //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (6),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("probs"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("probs_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_probs_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_6_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_6_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_probs_inst_dpi_control_done_writes_conduit),                    //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_probs_inst_dpi_control_done_reads_conduit),                     //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_6_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_6_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_probs_inst_m0_writedata),                                       //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_probs_inst_m0_burstcount),                                      //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdata),                                        //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_probs_inst_m0_address),                                         //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_probs_inst_m0_waitrequest),                                     //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_probs_inst_m0_write),                                           //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_probs_inst_m0_read),                                            //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_probs_inst_m0_byteenable),                                      //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdatavalid)                                    //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (5),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("w_conv1"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("w_conv1_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_w_conv1_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_7_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_7_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_w_conv1_inst_dpi_control_done_writes_conduit),                  //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_w_conv1_inst_dpi_control_done_reads_conduit),                   //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_7_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_7_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_writedata),                                     //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_burstcount),                                    //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdata),                                      //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_address),                                       //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_waitrequest),                                   //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_write),                                         //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_read),                                          //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_byteenable),                                    //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdatavalid)                                  //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (14),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("w_conv2"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("w_conv2_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_w_conv2_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_8_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_8_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_w_conv2_inst_dpi_control_done_writes_conduit),                  //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_w_conv2_inst_dpi_control_done_reads_conduit),                   //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_8_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_8_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_writedata),                                     //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_burstcount),                                    //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdata),                                      //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_address),                                       //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_waitrequest),                                   //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_write),                                         //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_read),                                          //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_byteenable),                                    //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdatavalid)                                  //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (18),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("w_fc1"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("w_fc1_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_w_fc1_inst (
		.clock              (clock_reset_inst_clock_clk),                                                             //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                           //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_9_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_9_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_w_fc1_inst_dpi_control_done_writes_conduit),                    //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_w_fc1_inst_dpi_control_done_reads_conduit),                     //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_9_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_9_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                       // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                       //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_writedata),                                       //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_burstcount),                                      //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdata),                                        //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_address),                                         //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_waitrequest),                                     //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_write),                                           //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_read),                                            //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_byteenable),                                      //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdatavalid)                                    //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (16),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("w_fc2"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("w_fc2_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_w_fc2_inst (
		.clock              (clock_reset_inst_clock_clk),                                                              //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                            //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_10_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_10_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_w_fc2_inst_dpi_control_done_writes_conduit),                     //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_w_fc2_inst_dpi_control_done_reads_conduit),                      //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_10_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_10_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                        // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                        //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_writedata),                                        //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_burstcount),                                       //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdata),                                         //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_address),                                          //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_waitrequest),                                      //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_write),                                            //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_read),                                             //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_byteenable),                                       //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdatavalid)                                     //                               .readdatavalid
	);

	hls_sim_mm_host_dpi_bfm #(
		.AV_ADDRESS_W                         (12),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("pred"),
		.COMPONENT_HAS_AGENT_RETURN           (0),
		.COMPONENT_AGENT_WRITE_INTERFACE_NAME ("w_fc3"),
		.COMPONENT_AGENT_READ_INTERFACE_NAME  ("w_fc3_avs_readback"),
		.COMPONENT_CRA_AGENT                  (0),
		.NUM_AGENT_MEMORIES                   (0)
	) mm_host_dpi_bfm_pred_avs_w_fc3_inst (
		.clock              (clock_reset_inst_clock_clk),                                                              //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                            //                          reset.reset_n
		.do_bind            (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_11_conduit),           //               dpi_control_bind.conduit
		.enable             (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_11_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_host_dpi_bfm_pred_avs_w_fc3_inst_dpi_control_done_writes_conduit),                     //        dpi_control_done_writes.conduit
		.done_reads         (mm_host_dpi_bfm_pred_avs_w_fc3_inst_dpi_control_done_reads_conduit),                      //         dpi_control_done_reads.conduit
		.component_started  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_11_conduit), //  dpi_control_component_started.conduit
		.component_done     (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_11_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (),                                                                                        // cra_control_done_writes_to_cra.conduit
		.agent_busy_out     (),                                                                                        //                 agent_busy_out.conduit
		.avm_writedata      (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_writedata),                                        //                             m0.writedata
		.avm_burstcount     (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_burstcount),                                       //                               .burstcount
		.avm_readdata       (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdata),                                         //                               .readdata
		.avm_address        (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_address),                                          //                               .address
		.avm_waitrequest    (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_waitrequest),                                      //                               .waitrequest
		.avm_write          (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_write),                                            //                               .write
		.avm_read           (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_read),                                             //                               .read
		.avm_byteenable     (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_byteenable),                                       //                               .byteenable
		.avm_readdatavalid  (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdatavalid)                                     //                               .readdatavalid
	);

	tb_pred_component_dpi_controller_agent_done_concatenate_inst pred_component_dpi_controller_agent_done_concatenate_inst (
		.out_conduit   (pred_component_dpi_controller_agent_done_concatenate_inst_out_conduit_conduit), //   out_conduit.conduit
		.in_conduit_0  (mm_host_dpi_bfm_pred_avs_b_conv1_inst_dpi_control_done_reads_conduit),          //  in_conduit_0.conduit
		.in_conduit_1  (mm_host_dpi_bfm_pred_avs_b_conv2_inst_dpi_control_done_reads_conduit),          //  in_conduit_1.conduit
		.in_conduit_2  (mm_host_dpi_bfm_pred_avs_b_fc1_inst_dpi_control_done_reads_conduit),            //  in_conduit_2.conduit
		.in_conduit_3  (mm_host_dpi_bfm_pred_avs_b_fc2_inst_dpi_control_done_reads_conduit),            //  in_conduit_3.conduit
		.in_conduit_4  (mm_host_dpi_bfm_pred_avs_b_fc3_inst_dpi_control_done_reads_conduit),            //  in_conduit_4.conduit
		.in_conduit_5  (mm_host_dpi_bfm_pred_avs_image_inst_dpi_control_done_reads_conduit),            //  in_conduit_5.conduit
		.in_conduit_6  (mm_host_dpi_bfm_pred_avs_probs_inst_dpi_control_done_reads_conduit),            //  in_conduit_6.conduit
		.in_conduit_7  (mm_host_dpi_bfm_pred_avs_w_conv1_inst_dpi_control_done_reads_conduit),          //  in_conduit_7.conduit
		.in_conduit_8  (mm_host_dpi_bfm_pred_avs_w_conv2_inst_dpi_control_done_reads_conduit),          //  in_conduit_8.conduit
		.in_conduit_9  (mm_host_dpi_bfm_pred_avs_w_fc1_inst_dpi_control_done_reads_conduit),            //  in_conduit_9.conduit
		.in_conduit_10 (mm_host_dpi_bfm_pred_avs_w_fc2_inst_dpi_control_done_reads_conduit),            // in_conduit_10.conduit
		.in_conduit_11 (mm_host_dpi_bfm_pred_avs_w_fc3_inst_dpi_control_done_reads_conduit)             // in_conduit_11.conduit
	);

	tb_pred_component_dpi_controller_agent_readback_fanout_inst pred_component_dpi_controller_agent_readback_fanout_inst (
		.in_conduit     (component_dpi_controller_pred_inst_readback_from_agents_conduit),                 //     in_conduit.conduit
		.out_conduit_0  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_0_conduit),  //  out_conduit_0.conduit
		.out_conduit_1  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_1_conduit),  //  out_conduit_1.conduit
		.out_conduit_2  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_2_conduit),  //  out_conduit_2.conduit
		.out_conduit_3  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_3_conduit),  //  out_conduit_3.conduit
		.out_conduit_4  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_4_conduit),  //  out_conduit_4.conduit
		.out_conduit_5  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_5_conduit),  //  out_conduit_5.conduit
		.out_conduit_6  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_6_conduit),  //  out_conduit_6.conduit
		.out_conduit_7  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_7_conduit),  //  out_conduit_7.conduit
		.out_conduit_8  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_8_conduit),  //  out_conduit_8.conduit
		.out_conduit_9  (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_9_conduit),  //  out_conduit_9.conduit
		.out_conduit_10 (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_10_conduit), // out_conduit_10.conduit
		.out_conduit_11 (pred_component_dpi_controller_agent_readback_fanout_inst_out_conduit_11_conduit)  // out_conduit_11.conduit
	);

	tb_pred_component_dpi_controller_agent_done_concatenate_inst pred_component_dpi_controller_agent_ready_concatenate_inst (
		.out_conduit   (pred_component_dpi_controller_agent_ready_concatenate_inst_out_conduit_conduit), //   out_conduit.conduit
		.in_conduit_0  (mm_host_dpi_bfm_pred_avs_b_conv1_inst_dpi_control_done_writes_conduit),          //  in_conduit_0.conduit
		.in_conduit_1  (mm_host_dpi_bfm_pred_avs_b_conv2_inst_dpi_control_done_writes_conduit),          //  in_conduit_1.conduit
		.in_conduit_2  (mm_host_dpi_bfm_pred_avs_b_fc1_inst_dpi_control_done_writes_conduit),            //  in_conduit_2.conduit
		.in_conduit_3  (mm_host_dpi_bfm_pred_avs_b_fc2_inst_dpi_control_done_writes_conduit),            //  in_conduit_3.conduit
		.in_conduit_4  (mm_host_dpi_bfm_pred_avs_b_fc3_inst_dpi_control_done_writes_conduit),            //  in_conduit_4.conduit
		.in_conduit_5  (mm_host_dpi_bfm_pred_avs_image_inst_dpi_control_done_writes_conduit),            //  in_conduit_5.conduit
		.in_conduit_6  (mm_host_dpi_bfm_pred_avs_probs_inst_dpi_control_done_writes_conduit),            //  in_conduit_6.conduit
		.in_conduit_7  (mm_host_dpi_bfm_pred_avs_w_conv1_inst_dpi_control_done_writes_conduit),          //  in_conduit_7.conduit
		.in_conduit_8  (mm_host_dpi_bfm_pred_avs_w_conv2_inst_dpi_control_done_writes_conduit),          //  in_conduit_8.conduit
		.in_conduit_9  (mm_host_dpi_bfm_pred_avs_w_fc1_inst_dpi_control_done_writes_conduit),            //  in_conduit_9.conduit
		.in_conduit_10 (mm_host_dpi_bfm_pred_avs_w_fc2_inst_dpi_control_done_writes_conduit),            // in_conduit_10.conduit
		.in_conduit_11 (mm_host_dpi_bfm_pred_avs_w_fc3_inst_dpi_control_done_writes_conduit)             // in_conduit_11.conduit
	);

	tb_pred_component_dpi_controller_agent_readback_fanout_inst pred_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit     (component_dpi_controller_pred_inst_dpi_control_bind_conduit),                   //     in_conduit.conduit
		.out_conduit_0  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),  //  out_conduit_0.conduit
		.out_conduit_1  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),  //  out_conduit_1.conduit
		.out_conduit_2  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),  //  out_conduit_2.conduit
		.out_conduit_3  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),  //  out_conduit_3.conduit
		.out_conduit_4  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),  //  out_conduit_4.conduit
		.out_conduit_5  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_5_conduit),  //  out_conduit_5.conduit
		.out_conduit_6  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_6_conduit),  //  out_conduit_6.conduit
		.out_conduit_7  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_7_conduit),  //  out_conduit_7.conduit
		.out_conduit_8  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_8_conduit),  //  out_conduit_8.conduit
		.out_conduit_9  (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_9_conduit),  //  out_conduit_9.conduit
		.out_conduit_10 (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_10_conduit), // out_conduit_10.conduit
		.out_conduit_11 (pred_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_11_conduit)  // out_conduit_11.conduit
	);

	tb_pred_component_dpi_controller_agent_readback_fanout_inst pred_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit     (component_dpi_controller_pred_inst_dpi_control_enable_conduit),                   //     in_conduit.conduit
		.out_conduit_0  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),  //  out_conduit_0.conduit
		.out_conduit_1  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),  //  out_conduit_1.conduit
		.out_conduit_2  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),  //  out_conduit_2.conduit
		.out_conduit_3  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),  //  out_conduit_3.conduit
		.out_conduit_4  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),  //  out_conduit_4.conduit
		.out_conduit_5  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_5_conduit),  //  out_conduit_5.conduit
		.out_conduit_6  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_6_conduit),  //  out_conduit_6.conduit
		.out_conduit_7  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_7_conduit),  //  out_conduit_7.conduit
		.out_conduit_8  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_8_conduit),  //  out_conduit_8.conduit
		.out_conduit_9  (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_9_conduit),  //  out_conduit_9.conduit
		.out_conduit_10 (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_10_conduit), // out_conduit_10.conduit
		.out_conduit_11 (pred_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_11_conduit)  // out_conduit_11.conduit
	);

	tb_pred_component_dpi_controller_agent_readback_fanout_inst pred_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit     (component_dpi_controller_pred_inst_read_implicit_streams_conduit),                        //     in_conduit.conduit
		.out_conduit_0  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit),  //  out_conduit_0.conduit
		.out_conduit_1  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit),  //  out_conduit_1.conduit
		.out_conduit_2  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit),  //  out_conduit_2.conduit
		.out_conduit_3  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit),  //  out_conduit_3.conduit
		.out_conduit_4  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_4_conduit),  //  out_conduit_4.conduit
		.out_conduit_5  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_5_conduit),  //  out_conduit_5.conduit
		.out_conduit_6  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_6_conduit),  //  out_conduit_6.conduit
		.out_conduit_7  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_7_conduit),  //  out_conduit_7.conduit
		.out_conduit_8  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_8_conduit),  //  out_conduit_8.conduit
		.out_conduit_9  (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_9_conduit),  //  out_conduit_9.conduit
		.out_conduit_10 (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_10_conduit), // out_conduit_10.conduit
		.out_conduit_11 (pred_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_11_conduit)  // out_conduit_11.conduit
	);

	tb_pred_inst pred_inst (
		.avs_b_conv1_read       (mm_interconnect_0_pred_inst_avs_b_conv1_read),              // avs_b_conv1.read
		.avs_b_conv1_readdata   (mm_interconnect_0_pred_inst_avs_b_conv1_readdata),          //            .readdata
		.avs_b_conv1_write      (mm_interconnect_0_pred_inst_avs_b_conv1_write),             //            .write
		.avs_b_conv1_writedata  (mm_interconnect_0_pred_inst_avs_b_conv1_writedata),         //            .writedata
		.avs_b_conv1_address    (mm_interconnect_0_pred_inst_avs_b_conv1_address),           //            .address
		.avs_b_conv1_byteenable (mm_interconnect_0_pred_inst_avs_b_conv1_byteenable),        //            .byteenable
		.avs_b_conv2_read       (mm_interconnect_1_pred_inst_avs_b_conv2_read),              // avs_b_conv2.read
		.avs_b_conv2_readdata   (mm_interconnect_1_pred_inst_avs_b_conv2_readdata),          //            .readdata
		.avs_b_conv2_write      (mm_interconnect_1_pred_inst_avs_b_conv2_write),             //            .write
		.avs_b_conv2_writedata  (mm_interconnect_1_pred_inst_avs_b_conv2_writedata),         //            .writedata
		.avs_b_conv2_address    (mm_interconnect_1_pred_inst_avs_b_conv2_address),           //            .address
		.avs_b_conv2_byteenable (mm_interconnect_1_pred_inst_avs_b_conv2_byteenable),        //            .byteenable
		.avs_b_fc1_read         (mm_interconnect_2_pred_inst_avs_b_fc1_read),                //   avs_b_fc1.read
		.avs_b_fc1_readdata     (mm_interconnect_2_pred_inst_avs_b_fc1_readdata),            //            .readdata
		.avs_b_fc1_write        (mm_interconnect_2_pred_inst_avs_b_fc1_write),               //            .write
		.avs_b_fc1_writedata    (mm_interconnect_2_pred_inst_avs_b_fc1_writedata),           //            .writedata
		.avs_b_fc1_address      (mm_interconnect_2_pred_inst_avs_b_fc1_address),             //            .address
		.avs_b_fc1_byteenable   (mm_interconnect_2_pred_inst_avs_b_fc1_byteenable),          //            .byteenable
		.avs_b_fc2_read         (mm_interconnect_3_pred_inst_avs_b_fc2_read),                //   avs_b_fc2.read
		.avs_b_fc2_readdata     (mm_interconnect_3_pred_inst_avs_b_fc2_readdata),            //            .readdata
		.avs_b_fc2_write        (mm_interconnect_3_pred_inst_avs_b_fc2_write),               //            .write
		.avs_b_fc2_writedata    (mm_interconnect_3_pred_inst_avs_b_fc2_writedata),           //            .writedata
		.avs_b_fc2_address      (mm_interconnect_3_pred_inst_avs_b_fc2_address),             //            .address
		.avs_b_fc2_byteenable   (mm_interconnect_3_pred_inst_avs_b_fc2_byteenable),          //            .byteenable
		.avs_b_fc3_read         (mm_interconnect_4_pred_inst_avs_b_fc3_read),                //   avs_b_fc3.read
		.avs_b_fc3_readdata     (mm_interconnect_4_pred_inst_avs_b_fc3_readdata),            //            .readdata
		.avs_b_fc3_write        (mm_interconnect_4_pred_inst_avs_b_fc3_write),               //            .write
		.avs_b_fc3_writedata    (mm_interconnect_4_pred_inst_avs_b_fc3_writedata),           //            .writedata
		.avs_b_fc3_address      (mm_interconnect_4_pred_inst_avs_b_fc3_address),             //            .address
		.avs_b_fc3_byteenable   (mm_interconnect_4_pred_inst_avs_b_fc3_byteenable),          //            .byteenable
		.avs_image_read         (mm_interconnect_5_pred_inst_avs_image_read),                //   avs_image.read
		.avs_image_readdata     (mm_interconnect_5_pred_inst_avs_image_readdata),            //            .readdata
		.avs_image_write        (mm_interconnect_5_pred_inst_avs_image_write),               //            .write
		.avs_image_writedata    (mm_interconnect_5_pred_inst_avs_image_writedata),           //            .writedata
		.avs_image_address      (mm_interconnect_5_pred_inst_avs_image_address),             //            .address
		.avs_image_byteenable   (mm_interconnect_5_pred_inst_avs_image_byteenable),          //            .byteenable
		.avs_probs_read         (mm_interconnect_6_pred_inst_avs_probs_read),                //   avs_probs.read
		.avs_probs_readdata     (mm_interconnect_6_pred_inst_avs_probs_readdata),            //            .readdata
		.avs_probs_write        (mm_interconnect_6_pred_inst_avs_probs_write),               //            .write
		.avs_probs_writedata    (mm_interconnect_6_pred_inst_avs_probs_writedata),           //            .writedata
		.avs_probs_address      (mm_interconnect_6_pred_inst_avs_probs_address),             //            .address
		.avs_probs_byteenable   (mm_interconnect_6_pred_inst_avs_probs_byteenable),          //            .byteenable
		.avs_w_conv1_read       (mm_interconnect_7_pred_inst_avs_w_conv1_read),              // avs_w_conv1.read
		.avs_w_conv1_readdata   (mm_interconnect_7_pred_inst_avs_w_conv1_readdata),          //            .readdata
		.avs_w_conv1_write      (mm_interconnect_7_pred_inst_avs_w_conv1_write),             //            .write
		.avs_w_conv1_writedata  (mm_interconnect_7_pred_inst_avs_w_conv1_writedata),         //            .writedata
		.avs_w_conv1_address    (mm_interconnect_7_pred_inst_avs_w_conv1_address),           //            .address
		.avs_w_conv1_byteenable (mm_interconnect_7_pred_inst_avs_w_conv1_byteenable),        //            .byteenable
		.avs_w_conv2_read       (mm_interconnect_8_pred_inst_avs_w_conv2_read),              // avs_w_conv2.read
		.avs_w_conv2_readdata   (mm_interconnect_8_pred_inst_avs_w_conv2_readdata),          //            .readdata
		.avs_w_conv2_write      (mm_interconnect_8_pred_inst_avs_w_conv2_write),             //            .write
		.avs_w_conv2_writedata  (mm_interconnect_8_pred_inst_avs_w_conv2_writedata),         //            .writedata
		.avs_w_conv2_address    (mm_interconnect_8_pred_inst_avs_w_conv2_address),           //            .address
		.avs_w_conv2_byteenable (mm_interconnect_8_pred_inst_avs_w_conv2_byteenable),        //            .byteenable
		.avs_w_fc1_read         (mm_interconnect_9_pred_inst_avs_w_fc1_read),                //   avs_w_fc1.read
		.avs_w_fc1_readdata     (mm_interconnect_9_pred_inst_avs_w_fc1_readdata),            //            .readdata
		.avs_w_fc1_write        (mm_interconnect_9_pred_inst_avs_w_fc1_write),               //            .write
		.avs_w_fc1_writedata    (mm_interconnect_9_pred_inst_avs_w_fc1_writedata),           //            .writedata
		.avs_w_fc1_address      (mm_interconnect_9_pred_inst_avs_w_fc1_address),             //            .address
		.avs_w_fc1_byteenable   (mm_interconnect_9_pred_inst_avs_w_fc1_byteenable),          //            .byteenable
		.avs_w_fc2_read         (mm_interconnect_10_pred_inst_avs_w_fc2_read),               //   avs_w_fc2.read
		.avs_w_fc2_readdata     (mm_interconnect_10_pred_inst_avs_w_fc2_readdata),           //            .readdata
		.avs_w_fc2_write        (mm_interconnect_10_pred_inst_avs_w_fc2_write),              //            .write
		.avs_w_fc2_writedata    (mm_interconnect_10_pred_inst_avs_w_fc2_writedata),          //            .writedata
		.avs_w_fc2_address      (mm_interconnect_10_pred_inst_avs_w_fc2_address),            //            .address
		.avs_w_fc2_byteenable   (mm_interconnect_10_pred_inst_avs_w_fc2_byteenable),         //            .byteenable
		.avs_w_fc3_read         (mm_interconnect_11_pred_inst_avs_w_fc3_read),               //   avs_w_fc3.read
		.avs_w_fc3_readdata     (mm_interconnect_11_pred_inst_avs_w_fc3_readdata),           //            .readdata
		.avs_w_fc3_write        (mm_interconnect_11_pred_inst_avs_w_fc3_write),              //            .write
		.avs_w_fc3_writedata    (mm_interconnect_11_pred_inst_avs_w_fc3_writedata),          //            .writedata
		.avs_w_fc3_address      (mm_interconnect_11_pred_inst_avs_w_fc3_address),            //            .address
		.avs_w_fc3_byteenable   (mm_interconnect_11_pred_inst_avs_w_fc3_byteenable),         //            .byteenable
		.start                  (component_dpi_controller_pred_inst_component_call_valid),   //        call.valid
		.busy                   (pred_inst_call_stall),                                      //            .stall
		.clock                  (clock_reset_inst_clock_clk),                                //       clock.clk
		.resetn                 (clock_reset_inst_reset_reset),                              //       reset.reset_n
		.done                   (pred_inst_return_valid),                                    //      return.valid
		.stall                  (component_dpi_controller_pred_inst_component_return_stall)  //            .stall
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    // out_conduit_0.conduit
	);

	tb_mm_interconnect_0 mm_interconnect_0 (
		.clock_reset_inst_clock_clk                                              (clock_reset_inst_clock_clk),                             //                                            clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                          // mm_host_dpi_bfm_pred_avs_b_conv1_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_waitrequest),   //                                                                  .waitrequest
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_burstcount),    //                                                                  .burstcount
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_byteenable),    //                                                                  .byteenable
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_read),          //                                                                  .read
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdata),      //                                                                  .readdata
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_readdatavalid), //                                                                  .readdatavalid
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_write),         //                                                                  .write
		.mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_b_conv1_inst_m0_writedata),     //                                                                  .writedata
		.pred_inst_avs_b_conv1_address                                           (mm_interconnect_0_pred_inst_avs_b_conv1_address),        //                                             pred_inst_avs_b_conv1.address
		.pred_inst_avs_b_conv1_write                                             (mm_interconnect_0_pred_inst_avs_b_conv1_write),          //                                                                  .write
		.pred_inst_avs_b_conv1_read                                              (mm_interconnect_0_pred_inst_avs_b_conv1_read),           //                                                                  .read
		.pred_inst_avs_b_conv1_readdata                                          (mm_interconnect_0_pred_inst_avs_b_conv1_readdata),       //                                                                  .readdata
		.pred_inst_avs_b_conv1_writedata                                         (mm_interconnect_0_pred_inst_avs_b_conv1_writedata),      //                                                                  .writedata
		.pred_inst_avs_b_conv1_byteenable                                        (mm_interconnect_0_pred_inst_avs_b_conv1_byteenable)      //                                                                  .byteenable
	);

	tb_mm_interconnect_1 mm_interconnect_1 (
		.clock_reset_inst_clock_clk                                              (clock_reset_inst_clock_clk),                             //                                            clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                          // mm_host_dpi_bfm_pred_avs_b_conv2_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_waitrequest),   //                                                                  .waitrequest
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_burstcount),    //                                                                  .burstcount
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_byteenable),    //                                                                  .byteenable
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_read),          //                                                                  .read
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdata),      //                                                                  .readdata
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_readdatavalid), //                                                                  .readdatavalid
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_write),         //                                                                  .write
		.mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_b_conv2_inst_m0_writedata),     //                                                                  .writedata
		.pred_inst_avs_b_conv2_address                                           (mm_interconnect_1_pred_inst_avs_b_conv2_address),        //                                             pred_inst_avs_b_conv2.address
		.pred_inst_avs_b_conv2_write                                             (mm_interconnect_1_pred_inst_avs_b_conv2_write),          //                                                                  .write
		.pred_inst_avs_b_conv2_read                                              (mm_interconnect_1_pred_inst_avs_b_conv2_read),           //                                                                  .read
		.pred_inst_avs_b_conv2_readdata                                          (mm_interconnect_1_pred_inst_avs_b_conv2_readdata),       //                                                                  .readdata
		.pred_inst_avs_b_conv2_writedata                                         (mm_interconnect_1_pred_inst_avs_b_conv2_writedata),      //                                                                  .writedata
		.pred_inst_avs_b_conv2_byteenable                                        (mm_interconnect_1_pred_inst_avs_b_conv2_byteenable)      //                                                                  .byteenable
	);

	tb_mm_interconnect_2 mm_interconnect_2 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_b_fc1_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_b_fc1_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_b_fc1_address                                           (mm_interconnect_2_pred_inst_avs_b_fc1_address),        //                                             pred_inst_avs_b_fc1.address
		.pred_inst_avs_b_fc1_write                                             (mm_interconnect_2_pred_inst_avs_b_fc1_write),          //                                                                .write
		.pred_inst_avs_b_fc1_read                                              (mm_interconnect_2_pred_inst_avs_b_fc1_read),           //                                                                .read
		.pred_inst_avs_b_fc1_readdata                                          (mm_interconnect_2_pred_inst_avs_b_fc1_readdata),       //                                                                .readdata
		.pred_inst_avs_b_fc1_writedata                                         (mm_interconnect_2_pred_inst_avs_b_fc1_writedata),      //                                                                .writedata
		.pred_inst_avs_b_fc1_byteenable                                        (mm_interconnect_2_pred_inst_avs_b_fc1_byteenable)      //                                                                .byteenable
	);

	tb_mm_interconnect_3 mm_interconnect_3 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_b_fc2_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_b_fc2_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_b_fc2_address                                           (mm_interconnect_3_pred_inst_avs_b_fc2_address),        //                                             pred_inst_avs_b_fc2.address
		.pred_inst_avs_b_fc2_write                                             (mm_interconnect_3_pred_inst_avs_b_fc2_write),          //                                                                .write
		.pred_inst_avs_b_fc2_read                                              (mm_interconnect_3_pred_inst_avs_b_fc2_read),           //                                                                .read
		.pred_inst_avs_b_fc2_readdata                                          (mm_interconnect_3_pred_inst_avs_b_fc2_readdata),       //                                                                .readdata
		.pred_inst_avs_b_fc2_writedata                                         (mm_interconnect_3_pred_inst_avs_b_fc2_writedata),      //                                                                .writedata
		.pred_inst_avs_b_fc2_byteenable                                        (mm_interconnect_3_pred_inst_avs_b_fc2_byteenable)      //                                                                .byteenable
	);

	tb_mm_interconnect_4 mm_interconnect_4 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_b_fc3_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_b_fc3_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_b_fc3_address                                           (mm_interconnect_4_pred_inst_avs_b_fc3_address),        //                                             pred_inst_avs_b_fc3.address
		.pred_inst_avs_b_fc3_write                                             (mm_interconnect_4_pred_inst_avs_b_fc3_write),          //                                                                .write
		.pred_inst_avs_b_fc3_read                                              (mm_interconnect_4_pred_inst_avs_b_fc3_read),           //                                                                .read
		.pred_inst_avs_b_fc3_readdata                                          (mm_interconnect_4_pred_inst_avs_b_fc3_readdata),       //                                                                .readdata
		.pred_inst_avs_b_fc3_writedata                                         (mm_interconnect_4_pred_inst_avs_b_fc3_writedata),      //                                                                .writedata
		.pred_inst_avs_b_fc3_byteenable                                        (mm_interconnect_4_pred_inst_avs_b_fc3_byteenable)      //                                                                .byteenable
	);

	tb_mm_interconnect_5 mm_interconnect_5 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_image_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_image_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_image_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_image_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_image_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_image_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_image_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_image_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_image_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_image_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_image_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_image_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_image_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_image_address                                           (mm_interconnect_5_pred_inst_avs_image_address),        //                                             pred_inst_avs_image.address
		.pred_inst_avs_image_write                                             (mm_interconnect_5_pred_inst_avs_image_write),          //                                                                .write
		.pred_inst_avs_image_read                                              (mm_interconnect_5_pred_inst_avs_image_read),           //                                                                .read
		.pred_inst_avs_image_readdata                                          (mm_interconnect_5_pred_inst_avs_image_readdata),       //                                                                .readdata
		.pred_inst_avs_image_writedata                                         (mm_interconnect_5_pred_inst_avs_image_writedata),      //                                                                .writedata
		.pred_inst_avs_image_byteenable                                        (mm_interconnect_5_pred_inst_avs_image_byteenable)      //                                                                .byteenable
	);

	tb_mm_interconnect_6 mm_interconnect_6 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_probs_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_probs_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_probs_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_probs_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_probs_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_probs_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_probs_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_probs_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_probs_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_probs_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_probs_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_probs_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_probs_address                                           (mm_interconnect_6_pred_inst_avs_probs_address),        //                                             pred_inst_avs_probs.address
		.pred_inst_avs_probs_write                                             (mm_interconnect_6_pred_inst_avs_probs_write),          //                                                                .write
		.pred_inst_avs_probs_read                                              (mm_interconnect_6_pred_inst_avs_probs_read),           //                                                                .read
		.pred_inst_avs_probs_readdata                                          (mm_interconnect_6_pred_inst_avs_probs_readdata),       //                                                                .readdata
		.pred_inst_avs_probs_writedata                                         (mm_interconnect_6_pred_inst_avs_probs_writedata),      //                                                                .writedata
		.pred_inst_avs_probs_byteenable                                        (mm_interconnect_6_pred_inst_avs_probs_byteenable)      //                                                                .byteenable
	);

	tb_mm_interconnect_7 mm_interconnect_7 (
		.clock_reset_inst_clock_clk                                              (clock_reset_inst_clock_clk),                             //                                            clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                          // mm_host_dpi_bfm_pred_avs_w_conv1_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_waitrequest),   //                                                                  .waitrequest
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_burstcount),    //                                                                  .burstcount
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_byteenable),    //                                                                  .byteenable
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_read),          //                                                                  .read
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdata),      //                                                                  .readdata
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_readdatavalid), //                                                                  .readdatavalid
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_write),         //                                                                  .write
		.mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_w_conv1_inst_m0_writedata),     //                                                                  .writedata
		.pred_inst_avs_w_conv1_address                                           (mm_interconnect_7_pred_inst_avs_w_conv1_address),        //                                             pred_inst_avs_w_conv1.address
		.pred_inst_avs_w_conv1_write                                             (mm_interconnect_7_pred_inst_avs_w_conv1_write),          //                                                                  .write
		.pred_inst_avs_w_conv1_read                                              (mm_interconnect_7_pred_inst_avs_w_conv1_read),           //                                                                  .read
		.pred_inst_avs_w_conv1_readdata                                          (mm_interconnect_7_pred_inst_avs_w_conv1_readdata),       //                                                                  .readdata
		.pred_inst_avs_w_conv1_writedata                                         (mm_interconnect_7_pred_inst_avs_w_conv1_writedata),      //                                                                  .writedata
		.pred_inst_avs_w_conv1_byteenable                                        (mm_interconnect_7_pred_inst_avs_w_conv1_byteenable)      //                                                                  .byteenable
	);

	tb_mm_interconnect_8 mm_interconnect_8 (
		.clock_reset_inst_clock_clk                                              (clock_reset_inst_clock_clk),                             //                                            clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                          // mm_host_dpi_bfm_pred_avs_w_conv2_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_waitrequest),   //                                                                  .waitrequest
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_burstcount),    //                                                                  .burstcount
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_byteenable),    //                                                                  .byteenable
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_read),          //                                                                  .read
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdata),      //                                                                  .readdata
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_readdatavalid), //                                                                  .readdatavalid
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_write),         //                                                                  .write
		.mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_w_conv2_inst_m0_writedata),     //                                                                  .writedata
		.pred_inst_avs_w_conv2_address                                           (mm_interconnect_8_pred_inst_avs_w_conv2_address),        //                                             pred_inst_avs_w_conv2.address
		.pred_inst_avs_w_conv2_write                                             (mm_interconnect_8_pred_inst_avs_w_conv2_write),          //                                                                  .write
		.pred_inst_avs_w_conv2_read                                              (mm_interconnect_8_pred_inst_avs_w_conv2_read),           //                                                                  .read
		.pred_inst_avs_w_conv2_readdata                                          (mm_interconnect_8_pred_inst_avs_w_conv2_readdata),       //                                                                  .readdata
		.pred_inst_avs_w_conv2_writedata                                         (mm_interconnect_8_pred_inst_avs_w_conv2_writedata),      //                                                                  .writedata
		.pred_inst_avs_w_conv2_byteenable                                        (mm_interconnect_8_pred_inst_avs_w_conv2_byteenable)      //                                                                  .byteenable
	);

	tb_mm_interconnect_9 mm_interconnect_9 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_w_fc1_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_w_fc1_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_w_fc1_address                                           (mm_interconnect_9_pred_inst_avs_w_fc1_address),        //                                             pred_inst_avs_w_fc1.address
		.pred_inst_avs_w_fc1_write                                             (mm_interconnect_9_pred_inst_avs_w_fc1_write),          //                                                                .write
		.pred_inst_avs_w_fc1_read                                              (mm_interconnect_9_pred_inst_avs_w_fc1_read),           //                                                                .read
		.pred_inst_avs_w_fc1_readdata                                          (mm_interconnect_9_pred_inst_avs_w_fc1_readdata),       //                                                                .readdata
		.pred_inst_avs_w_fc1_writedata                                         (mm_interconnect_9_pred_inst_avs_w_fc1_writedata),      //                                                                .writedata
		.pred_inst_avs_w_fc1_byteenable                                        (mm_interconnect_9_pred_inst_avs_w_fc1_byteenable)      //                                                                .byteenable
	);

	tb_mm_interconnect_10 mm_interconnect_10 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_w_fc2_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_w_fc2_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_w_fc2_address                                           (mm_interconnect_10_pred_inst_avs_w_fc2_address),       //                                             pred_inst_avs_w_fc2.address
		.pred_inst_avs_w_fc2_write                                             (mm_interconnect_10_pred_inst_avs_w_fc2_write),         //                                                                .write
		.pred_inst_avs_w_fc2_read                                              (mm_interconnect_10_pred_inst_avs_w_fc2_read),          //                                                                .read
		.pred_inst_avs_w_fc2_readdata                                          (mm_interconnect_10_pred_inst_avs_w_fc2_readdata),      //                                                                .readdata
		.pred_inst_avs_w_fc2_writedata                                         (mm_interconnect_10_pred_inst_avs_w_fc2_writedata),     //                                                                .writedata
		.pred_inst_avs_w_fc2_byteenable                                        (mm_interconnect_10_pred_inst_avs_w_fc2_byteenable)     //                                                                .byteenable
	);

	tb_mm_interconnect_11 mm_interconnect_11 (
		.clock_reset_inst_clock_clk                                            (clock_reset_inst_clock_clk),                           //                                          clock_reset_inst_clock.clk
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                        // mm_host_dpi_bfm_pred_avs_w_fc3_inst_reset_reset_bridge_in_reset.reset
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_address                        (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_address),       //                          mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0.address
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_waitrequest                    (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_waitrequest),   //                                                                .waitrequest
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_burstcount                     (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_burstcount),    //                                                                .burstcount
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_byteenable                     (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_byteenable),    //                                                                .byteenable
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_read                           (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_read),          //                                                                .read
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdata                       (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdata),      //                                                                .readdata
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdatavalid                  (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_readdatavalid), //                                                                .readdatavalid
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_write                          (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_write),         //                                                                .write
		.mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_writedata                      (mm_host_dpi_bfm_pred_avs_w_fc3_inst_m0_writedata),     //                                                                .writedata
		.pred_inst_avs_w_fc3_address                                           (mm_interconnect_11_pred_inst_avs_w_fc3_address),       //                                             pred_inst_avs_w_fc3.address
		.pred_inst_avs_w_fc3_write                                             (mm_interconnect_11_pred_inst_avs_w_fc3_write),         //                                                                .write
		.pred_inst_avs_w_fc3_read                                              (mm_interconnect_11_pred_inst_avs_w_fc3_read),          //                                                                .read
		.pred_inst_avs_w_fc3_readdata                                          (mm_interconnect_11_pred_inst_avs_w_fc3_readdata),      //                                                                .readdata
		.pred_inst_avs_w_fc3_writedata                                         (mm_interconnect_11_pred_inst_avs_w_fc3_writedata),     //                                                                .writedata
		.pred_inst_avs_w_fc3_byteenable                                        (mm_interconnect_11_pred_inst_avs_w_fc3_byteenable)     //                                                                .byteenable
	);

	tb_irq_mapper irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                           //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                        // clk_reset.reset
		.sender_irq (component_dpi_controller_pred_inst_component_irq_irq)  //    sender.irq
	);

endmodule
