// tb.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module tb (
	);

	wire         clock_reset_inst_clock_clk;                                                            // clock_reset_inst:clock -> [component_dpi_controller_dut_inst:clock, dut_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock, stream_source_dpi_bfm_dut_x_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                          // clock_reset_inst:clock2x -> [component_dpi_controller_dut_inst:clock2x, main_dpi_controller_inst:clock2x, stream_source_dpi_bfm_dut_x_inst:clock2x]
	wire         component_dpi_controller_dut_inst_component_call_valid;                                // component_dpi_controller_dut_inst:start -> dut_inst:start
	wire         dut_inst_call_stall;                                                                   // dut_inst:busy -> component_dpi_controller_dut_inst:busy
	wire         component_dpi_controller_dut_inst_component_done_conduit;                              // component_dpi_controller_dut_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire   [0:0] main_dpi_controller_inst_component_enabled_conduit;                                    // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_dut_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_dut_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         component_dpi_controller_dut_inst_dpi_control_bind_conduit;                            // component_dpi_controller_dut_inst:bind_interfaces -> dut_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_dut_inst_dpi_control_enable_conduit;                          // component_dpi_controller_dut_inst:enable_interfaces -> dut_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         concatenate_component_done_inst_out_conduit_conduit;                                   // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire         concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                 // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire         split_component_start_inst_out_conduit_0_conduit;                                      // split_component_start_inst:out_conduit_0 -> component_dpi_controller_dut_inst:component_enabled
	wire         dut_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // dut_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_dut_x_inst:do_bind
	wire         dut_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // dut_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_dut_x_inst:enable
	wire         dut_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // dut_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_dut_x_inst:source_ready
	wire         component_dpi_controller_dut_inst_read_implicit_streams_conduit;                       // component_dpi_controller_dut_inst:read_implicit_streams -> dut_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                           // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         dut_inst_return_valid;                                                                 // dut_inst:done -> component_dpi_controller_dut_inst:done
	wire         component_dpi_controller_dut_inst_component_return_stall;                              // component_dpi_controller_dut_inst:stall -> dut_inst:stall
	wire  [15:0] dut_inst_returndata_data;                                                              // dut_inst:returndata -> component_dpi_controller_dut_inst:returndata
	wire  [15:0] stream_source_dpi_bfm_dut_x_inst_source_data_data;                                     // stream_source_dpi_bfm_dut_x_inst:source_data -> dut_inst:x
	wire         clock_reset_inst_reset_reset;                                                          // clock_reset_inst:resetn -> [component_dpi_controller_dut_inst:resetn, dut_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn, stream_source_dpi_bfm_dut_x_inst:resetn]
	wire         component_dpi_controller_dut_inst_component_irq_irq;                                   // irq_mapper:sender_irq -> component_dpi_controller_dut_inst:done_irq

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("dut"),
		.COMPONENT_MANGLED_NAME       ("\\3fdut@@YA\\3fAV\\3f$ac_fixed@$0BA@$07$00$0A@$0A@@@V1@@Z"),
		.RETURN_DATAWIDTH             (16),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_dut_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                 //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                               //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                               //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_dut_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_dut_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                           //                component_enabled.conduit
		.component_done                   (component_dpi_controller_dut_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_dut_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                           //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_dut_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                           //             readback_from_agents.conduit
		.start                            (component_dpi_controller_dut_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (dut_inst_call_stall),                                                        //                                 .stall
		.done                             (dut_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_dut_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_dut_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       (dut_inst_returndata_data)                                                    //                       returndata.data
	);

	tb_concatenate_component_done_inst concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),      //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_dut_inst_component_done_conduit)  // in_conduit_0.conduit
	);

	tb_concatenate_component_done_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),      //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_dut_inst_component_wait_for_stream_writes_conduit)  // in_conduit_0.conduit
	);

	tb_dut_component_dpi_controller_bind_conduit_fanout_inst dut_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_dut_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (dut_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit)  // out_conduit_0.conduit
	);

	tb_dut_component_dpi_controller_bind_conduit_fanout_inst dut_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_dut_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (dut_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit)  // out_conduit_0.conduit
	);

	tb_dut_component_dpi_controller_bind_conduit_fanout_inst dut_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_dut_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (dut_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit)  // out_conduit_0.conduit
	);

	tb_dut_inst dut_inst (
		.start      (component_dpi_controller_dut_inst_component_call_valid),   //       call.valid
		.busy       (dut_inst_call_stall),                                      //           .stall
		.clock      (clock_reset_inst_clock_clk),                               //      clock.clk
		.resetn     (clock_reset_inst_reset_reset),                             //      reset.reset_n
		.done       (dut_inst_return_valid),                                    //     return.valid
		.stall      (component_dpi_controller_dut_inst_component_return_stall), //           .stall
		.returndata (dut_inst_returndata_data),                                 // returndata.data
		.x          (stream_source_dpi_bfm_dut_x_inst_source_data_data)         //          x.data
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS      (1),
		.COMPONENT_NAMES_STR ("dut")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    // out_conduit_0.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("dut"),
		.INTERFACE_NAME                  ("x"),
		.STREAM_DATAWIDTH                (16),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_dut_x_inst (
		.clock        (clock_reset_inst_clock_clk),                                                            //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                          //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                          //            clock2x.clk
		.do_bind      (dut_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),           //   dpi_control_bind.conduit
		.enable       (dut_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_dut_x_inst_source_data_data),                                     //        source_data.data
		.source_ready (dut_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                       //             source.conduit
	);

	tb_irq_mapper irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                          //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                       // clk_reset.reset
		.sender_irq (component_dpi_controller_dut_inst_component_irq_irq)  //    sender.irq
	);

endmodule
