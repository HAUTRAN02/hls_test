// tb_dut_inst.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module tb_dut_inst (
		input  wire        start,      //       call.valid
		output wire        busy,       //           .stall
		input  wire        clock,      //      clock.clk
		input  wire        resetn,     //      reset.reset_n
		output wire        done,       //     return.valid
		input  wire        stall,      //           .stall
		output wire [15:0] returndata, // returndata.data
		input  wire [15:0] x           //          x.data
	);

	dut_internal dut_internal_inst (
		.clock      (clock),      //      clock.clk
		.resetn     (resetn),     //      reset.reset_n
		.start      (start),      //       call.valid
		.busy       (busy),       //           .stall
		.done       (done),       //     return.valid
		.stall      (stall),      //           .stall
		.returndata (returndata), // returndata.data
		.x          (x)           //          x.data
	);

endmodule
