// tb_pred_inst.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module tb_pred_inst (
		input  wire        avs_b_conv1_read,       // avs_b_conv1.read
		output wire [31:0] avs_b_conv1_readdata,   //            .readdata
		input  wire        avs_b_conv1_write,      //            .write
		input  wire [31:0] avs_b_conv1_writedata,  //            .writedata
		input  wire [2:0]  avs_b_conv1_address,    //            .address
		input  wire [3:0]  avs_b_conv1_byteenable, //            .byteenable
		input  wire        avs_b_conv2_read,       // avs_b_conv2.read
		output wire [31:0] avs_b_conv2_readdata,   //            .readdata
		input  wire        avs_b_conv2_write,      //            .write
		input  wire [31:0] avs_b_conv2_writedata,  //            .writedata
		input  wire [3:0]  avs_b_conv2_address,    //            .address
		input  wire [3:0]  avs_b_conv2_byteenable, //            .byteenable
		input  wire        avs_b_fc1_read,         //   avs_b_fc1.read
		output wire [31:0] avs_b_fc1_readdata,     //            .readdata
		input  wire        avs_b_fc1_write,        //            .write
		input  wire [31:0] avs_b_fc1_writedata,    //            .writedata
		input  wire [6:0]  avs_b_fc1_address,      //            .address
		input  wire [3:0]  avs_b_fc1_byteenable,   //            .byteenable
		input  wire        avs_b_fc2_read,         //   avs_b_fc2.read
		output wire [31:0] avs_b_fc2_readdata,     //            .readdata
		input  wire        avs_b_fc2_write,        //            .write
		input  wire [31:0] avs_b_fc2_writedata,    //            .writedata
		input  wire [6:0]  avs_b_fc2_address,      //            .address
		input  wire [3:0]  avs_b_fc2_byteenable,   //            .byteenable
		input  wire        avs_b_fc3_read,         //   avs_b_fc3.read
		output wire [31:0] avs_b_fc3_readdata,     //            .readdata
		input  wire        avs_b_fc3_write,        //            .write
		input  wire [31:0] avs_b_fc3_writedata,    //            .writedata
		input  wire [3:0]  avs_b_fc3_address,      //            .address
		input  wire [3:0]  avs_b_fc3_byteenable,   //            .byteenable
		input  wire        avs_image_read,         //   avs_image.read
		output wire [31:0] avs_image_readdata,     //            .readdata
		input  wire        avs_image_write,        //            .write
		input  wire [31:0] avs_image_writedata,    //            .writedata
		input  wire [9:0]  avs_image_address,      //            .address
		input  wire [3:0]  avs_image_byteenable,   //            .byteenable
		input  wire        avs_probs_read,         //   avs_probs.read
		output wire [31:0] avs_probs_readdata,     //            .readdata
		input  wire        avs_probs_write,        //            .write
		input  wire [31:0] avs_probs_writedata,    //            .writedata
		input  wire [3:0]  avs_probs_address,      //            .address
		input  wire [3:0]  avs_probs_byteenable,   //            .byteenable
		input  wire        avs_w_conv1_read,       // avs_w_conv1.read
		output wire [31:0] avs_w_conv1_readdata,   //            .readdata
		input  wire        avs_w_conv1_write,      //            .write
		input  wire [31:0] avs_w_conv1_writedata,  //            .writedata
		input  wire [2:0]  avs_w_conv1_address,    //            .address
		input  wire [3:0]  avs_w_conv1_byteenable, //            .byteenable
		input  wire        avs_w_conv2_read,       // avs_w_conv2.read
		output wire [31:0] avs_w_conv2_readdata,   //            .readdata
		input  wire        avs_w_conv2_write,      //            .write
		input  wire [31:0] avs_w_conv2_writedata,  //            .writedata
		input  wire [11:0] avs_w_conv2_address,    //            .address
		input  wire [3:0]  avs_w_conv2_byteenable, //            .byteenable
		input  wire        avs_w_fc1_read,         //   avs_w_fc1.read
		output wire [31:0] avs_w_fc1_readdata,     //            .readdata
		input  wire        avs_w_fc1_write,        //            .write
		input  wire [31:0] avs_w_fc1_writedata,    //            .writedata
		input  wire [15:0] avs_w_fc1_address,      //            .address
		input  wire [3:0]  avs_w_fc1_byteenable,   //            .byteenable
		input  wire        avs_w_fc2_read,         //   avs_w_fc2.read
		output wire [31:0] avs_w_fc2_readdata,     //            .readdata
		input  wire        avs_w_fc2_write,        //            .write
		input  wire [31:0] avs_w_fc2_writedata,    //            .writedata
		input  wire [13:0] avs_w_fc2_address,      //            .address
		input  wire [3:0]  avs_w_fc2_byteenable,   //            .byteenable
		input  wire        avs_w_fc3_read,         //   avs_w_fc3.read
		output wire [31:0] avs_w_fc3_readdata,     //            .readdata
		input  wire        avs_w_fc3_write,        //            .write
		input  wire [31:0] avs_w_fc3_writedata,    //            .writedata
		input  wire [9:0]  avs_w_fc3_address,      //            .address
		input  wire [3:0]  avs_w_fc3_byteenable,   //            .byteenable
		input  wire        start,                  //        call.valid
		output wire        busy,                   //            .stall
		input  wire        clock,                  //       clock.clk
		input  wire        resetn,                 //       reset.reset_n
		output wire        done,                   //      return.valid
		input  wire        stall                   //            .stall
	);

	pred_internal pred_internal_inst (
		.clock                  (clock),                  //       clock.clk
		.resetn                 (resetn),                 //       reset.reset_n
		.start                  (start),                  //        call.valid
		.busy                   (busy),                   //            .stall
		.done                   (done),                   //      return.valid
		.stall                  (stall),                  //            .stall
		.avs_b_conv1_read       (avs_b_conv1_read),       // avs_b_conv1.read
		.avs_b_conv1_readdata   (avs_b_conv1_readdata),   //            .readdata
		.avs_b_conv1_write      (avs_b_conv1_write),      //            .write
		.avs_b_conv1_writedata  (avs_b_conv1_writedata),  //            .writedata
		.avs_b_conv1_address    (avs_b_conv1_address),    //            .address
		.avs_b_conv1_byteenable (avs_b_conv1_byteenable), //            .byteenable
		.avs_b_conv2_read       (avs_b_conv2_read),       // avs_b_conv2.read
		.avs_b_conv2_readdata   (avs_b_conv2_readdata),   //            .readdata
		.avs_b_conv2_write      (avs_b_conv2_write),      //            .write
		.avs_b_conv2_writedata  (avs_b_conv2_writedata),  //            .writedata
		.avs_b_conv2_address    (avs_b_conv2_address),    //            .address
		.avs_b_conv2_byteenable (avs_b_conv2_byteenable), //            .byteenable
		.avs_b_fc1_read         (avs_b_fc1_read),         //   avs_b_fc1.read
		.avs_b_fc1_readdata     (avs_b_fc1_readdata),     //            .readdata
		.avs_b_fc1_write        (avs_b_fc1_write),        //            .write
		.avs_b_fc1_writedata    (avs_b_fc1_writedata),    //            .writedata
		.avs_b_fc1_address      (avs_b_fc1_address),      //            .address
		.avs_b_fc1_byteenable   (avs_b_fc1_byteenable),   //            .byteenable
		.avs_b_fc2_read         (avs_b_fc2_read),         //   avs_b_fc2.read
		.avs_b_fc2_readdata     (avs_b_fc2_readdata),     //            .readdata
		.avs_b_fc2_write        (avs_b_fc2_write),        //            .write
		.avs_b_fc2_writedata    (avs_b_fc2_writedata),    //            .writedata
		.avs_b_fc2_address      (avs_b_fc2_address),      //            .address
		.avs_b_fc2_byteenable   (avs_b_fc2_byteenable),   //            .byteenable
		.avs_b_fc3_read         (avs_b_fc3_read),         //   avs_b_fc3.read
		.avs_b_fc3_readdata     (avs_b_fc3_readdata),     //            .readdata
		.avs_b_fc3_write        (avs_b_fc3_write),        //            .write
		.avs_b_fc3_writedata    (avs_b_fc3_writedata),    //            .writedata
		.avs_b_fc3_address      (avs_b_fc3_address),      //            .address
		.avs_b_fc3_byteenable   (avs_b_fc3_byteenable),   //            .byteenable
		.avs_image_read         (avs_image_read),         //   avs_image.read
		.avs_image_readdata     (avs_image_readdata),     //            .readdata
		.avs_image_write        (avs_image_write),        //            .write
		.avs_image_writedata    (avs_image_writedata),    //            .writedata
		.avs_image_address      (avs_image_address),      //            .address
		.avs_image_byteenable   (avs_image_byteenable),   //            .byteenable
		.avs_probs_read         (avs_probs_read),         //   avs_probs.read
		.avs_probs_readdata     (avs_probs_readdata),     //            .readdata
		.avs_probs_write        (avs_probs_write),        //            .write
		.avs_probs_writedata    (avs_probs_writedata),    //            .writedata
		.avs_probs_address      (avs_probs_address),      //            .address
		.avs_probs_byteenable   (avs_probs_byteenable),   //            .byteenable
		.avs_w_conv1_read       (avs_w_conv1_read),       // avs_w_conv1.read
		.avs_w_conv1_readdata   (avs_w_conv1_readdata),   //            .readdata
		.avs_w_conv1_write      (avs_w_conv1_write),      //            .write
		.avs_w_conv1_writedata  (avs_w_conv1_writedata),  //            .writedata
		.avs_w_conv1_address    (avs_w_conv1_address),    //            .address
		.avs_w_conv1_byteenable (avs_w_conv1_byteenable), //            .byteenable
		.avs_w_conv2_read       (avs_w_conv2_read),       // avs_w_conv2.read
		.avs_w_conv2_readdata   (avs_w_conv2_readdata),   //            .readdata
		.avs_w_conv2_write      (avs_w_conv2_write),      //            .write
		.avs_w_conv2_writedata  (avs_w_conv2_writedata),  //            .writedata
		.avs_w_conv2_address    (avs_w_conv2_address),    //            .address
		.avs_w_conv2_byteenable (avs_w_conv2_byteenable), //            .byteenable
		.avs_w_fc1_read         (avs_w_fc1_read),         //   avs_w_fc1.read
		.avs_w_fc1_readdata     (avs_w_fc1_readdata),     //            .readdata
		.avs_w_fc1_write        (avs_w_fc1_write),        //            .write
		.avs_w_fc1_writedata    (avs_w_fc1_writedata),    //            .writedata
		.avs_w_fc1_address      (avs_w_fc1_address),      //            .address
		.avs_w_fc1_byteenable   (avs_w_fc1_byteenable),   //            .byteenable
		.avs_w_fc2_read         (avs_w_fc2_read),         //   avs_w_fc2.read
		.avs_w_fc2_readdata     (avs_w_fc2_readdata),     //            .readdata
		.avs_w_fc2_write        (avs_w_fc2_write),        //            .write
		.avs_w_fc2_writedata    (avs_w_fc2_writedata),    //            .writedata
		.avs_w_fc2_address      (avs_w_fc2_address),      //            .address
		.avs_w_fc2_byteenable   (avs_w_fc2_byteenable),   //            .byteenable
		.avs_w_fc3_read         (avs_w_fc3_read),         //   avs_w_fc3.read
		.avs_w_fc3_readdata     (avs_w_fc3_readdata),     //            .readdata
		.avs_w_fc3_write        (avs_w_fc3_write),        //            .write
		.avs_w_fc3_writedata    (avs_w_fc3_writedata),    //            .writedata
		.avs_w_fc3_address      (avs_w_fc3_address),      //            .address
		.avs_w_fc3_byteenable   (avs_w_fc3_byteenable)    //            .byteenable
	);

endmodule
